module SPI_mnrch(
	input 				clk, rst_n,
	input 				wrt,
	input [15:0]		wt_data,
	input 				MISO,
	output 				SS_n,
	output 				SCLK,
	output 				MOSI,
	output 				done,
	output [15:0]		rd_data
);
	// SCLK counter and signals
	logic [4:0] SCLK_div;
	logic SCLK_fall, SCLK_rise;
	
	// bit counter
	logic [3:0] bit_cnt;
	logic done15;
	
	// 16-bit shift register
	logic [15:0] shft_reg;
	logic MISO_smpl;

	// SM outputs
	logic smpl, init, shift, rst_cnt, set_done, ld_SCLK;
	
	typedef enum reg [1:0] { IDLE, SKIP, WAIT15, DONE } state_t;
	state_t state, nxt_state;

	////////// SCLK datapath //////////
	// 5-bit SCLK counter (requires preset since SCLK normally high)
	always_ff @(posedge clk, negedge rst_n)
		if(!rst_n)
			SCLK_div <= 5'h10;
		else if(ld_SCLK)
			SCLK_div <= 5'h17;
		else if()
			SCLK_div <= SCLK_div + 1;
		
	// SS_n
	always @(posedge clk, negedge rst_n)
		if(!rst_n)
			SS_n <= 1;
		else if(done)
			SS_n <= 1;
		else if(init)
			SS_n <= 0;
		
	assign SCLK = SCLK_div[4];
	assign shift = &SCLK_div;
	
	// imminent fall/rise
	assign SCLK_fall = ~SCLK_ff1 & SCLK_ff2;
	assign SCLK_rise = SCLK_ff1 & ~SCLK_ff2;
	
	
	/////// bit counter datapath ///////
	always_ff @(posedge clk)
		if(init)
			bit_cnt <= 4'h0;
		else if(shift)
			bit_cnt <= bit_cnt + 1;
			
	assign done15 = &bit_cnt;
	
	////////// shift register /////////
	always_ff @(posedge clk, negedge rst_n)
		if(smpl)
			MISO_smpl <= MISO;

	always_ff @(posedge clk, negedge rst_n)
		if(!rst_n)
			shft_reg <= 16'hFFFF;
		else if(init)
			shft_reg <= wt_data;
		else if(shift)
			shft_reg <= {shft_reg[14:0],MISO_smpl};

	assign MOSI = shft_reg[15];
	
	////////// state machine //////////
	// state register
	always_ff @(posedge clk, negedge rst_n)
		if(!rst_n)
			state <= IDLE;
		else
			state <= nxt_state;
	
	// TODO: output and transition logic
	always_comb begin
		nxt_state = state;
		case(state)
		
		endcase
	end
	
	// SR flop for done
	always_ff @(posedge clk, negedge rst_n)
		if(!rst_n)
			done <= 0;
		else if(init)
			done <= 0;
		else if(set_done)
			done <= 1;
endmodule